Circuito 2 

I1 0 n1 DC 1
R1 n1 n2 90
R2 n2 n6 80 
R3 n2 n5 40
R4 n2 0 10
R5 n2 n4 20 
R6 n4 n5 20
R7 n5 0 50 
R8 n6 n7 90 
R9 n5 n6 70
I2 0 n7 Dc 1 
V1 n4 0 DC 10
.end 

