Baticircuito
R1 n3 n7 1000
R3 n3 n5 3000
R4 n3 n4 4000
I5 n4 n3 DC 0.005 
R5 n3 n2 3000
R6 n3 n2 1000
R7 n5 n7 4000
R8 n5 n4 1000
R9 n4 n6 5000
R11 n4 n2 3000
R12 n7 n8 2000
R10 n6 n8 4000
I1 n1 n6 DC 0.001
R13 n6 n2 4000
R14 n2 n1 3000
R2 n1 n8 2000
R15 n8 n10 1000
R16 n8 n11 2000
R17 n10 n11 2000
R18 n8 n9 3000
I2 n9 n11 DC 0.002
R19 n10 n18 5000
R20 n9 n10 1000
R21 n18 n14 2000
R22 n10 n17 4000
R23 n9 n17 5000
R24 n9 n1 4000
R25 n1 0 3000
R26 n17 0 4000
I3 n17 n12 DC 0.003
R27 n18 n13 3000
R28 n13 n14 4000
R29 n12 n15 3000
R30 n13 n15 1000
R31 n15 n14 5000
R32 n17 n16 3000
R33 n12 n16 4000
R34 n16 n14 5000
R35 n16 n14 3000
R36 n16 n15 2000
R37 n10 n12 2000
I4 n14 n15 DC 0.004
.end
